module HistogramDisplayer(
	input iClk,
	input iRst_n,
	input [15:0] X_Cont,
	input [15:0] Y_Cont, 
	output 
						)